LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

LIBRARY work;
USE work.PCK_CRC32_D4.ALL;
USE work.common.ALL;

ENTITY mac_snd IS
  PORT (
    E_TX_CLK : IN STD_LOGIC; -- Sender Clock.
    E_TX_EN : OUT STD_LOGIC; -- Sender Enable.
    E_TXD : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- Sent Data.
    E_TX_ER : OUT STD_LOGIC; -- Sent Data Error.
    el_data : IN data_t; -- Actual data.
    el_snd_en : IN STD_LOGIC -- User Start Send.
  );
END mac_snd;

ARCHITECTURE rtl OF mac_snd IS

  TYPE mem_t IS ARRAY(0 TO 14) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

  -- -- TO BE REMOVED
  -- SIGNAL mem : mem_t := (
  --   -- DST MAC Address
  --   x"00", x"e0", x"4c", x"6b", x"dc", x"98",

  --   -- FPGA MAC Address (Xilinx OUI)                                        --
  --   x"00", x"0a", x"35", x"00", x"00", x"00",

  --   -- EtherType Field: 0x0000                                              --
  --   x"08", x"00",

  --   -- Data Header                                                          --
  --   x"45"
  -- );

  --ATTRIBUTE RAM_STYLE : STRING;
  --ATTRIBUTE RAM_STYLE OF mem : SIGNAL IS "BLOCK";

  TYPE state_t IS (
    Idle, -- Wait for signal en.
    Preamble, -- 55 55 55 55 55 55 55 5
    StartOfFrame, -- d
    --EtherUpper, -- 6 Byte MAC address Upper nibble
    --EtherLower, -- 6 Byte MAC address Lower nibble
    EtherMACDST, -- 6 Byte MAC DST address
    EtherMACSRC, -- 6 Byte MAC SRC address
    EtherType, -- 0x0800
    IPVersion, -- 0x4
    IPIHL, -- 0x5
    IPDSCPECN, -- 0x00
    IPLength, -- ipLength
    IPID, -- 0x00
    IPFlagsFragment, -- 0x00
    IPTTL, -- 0x40
    IPProtocol, -- 0x11
    IPChecksum, -- Checksum
    IPAddrSRC, -- IPAddr SRC
    IPAddrDST, -- IPAddr DST
    -- UDPPortSRC, -- 2 byte UDP SRC
    -- UDPPortDST, -- 2 byte UDP DST
    -- UDPChecksum, -- Checksum,
    DNSMsg, -- 1472 Max bytes
    FrameCheck, -- CRC32
    InterframeGap -- Gap between two cosecutive frames (24 Bit).
  );

  TYPE snd_t IS RECORD
    s : state_t;
    d : data_t;
    crc : STD_LOGIC_VECTOR(31 DOWNTO 0); -- CRC32 latch.
    c : NATURAL RANGE 0 TO 367;
  END RECORD;

  SIGNAL s, sin : snd_t
    := snd_t'(
      s => Idle,
      d => (
        srcMAC => (OTHERS => '0'), dstMAC => (OTHERS => '0'),
        srcIP  => (OTHERS => '0'), dstIP => (OTHERS => '0'),
        ipHeaderLength => 0, ipLength => 0,
        srcPort => (OTHERS => '0'), dstPort => (OTHERS => '0'), dnsLength => 0
        --dns => (OTHERS => '0')
      ),
      crc => x"ffffffff",
      c => 0
    );

BEGIN

  snd_nsl : PROCESS (s, el_snd_en, el_data) -- mem
  BEGIN

    sin <= s;
    E_TX_EN <= '0';
    E_TXD <= x"0";
    E_TX_ER <= '0';

    CASE s.s IS
      WHEN Idle =>
        IF el_snd_en = '1' THEN
          sin.c <= 0;
          sin.s <= Preamble;
          sin.d <= el_data;
        END IF;

      -- Preamble, 15 5s (including nibble for start of frame)
      WHEN Preamble =>
        E_TXD <= x"5";
        E_TX_EN <= '1';
        IF s.c = 14 THEN
          sin.c <= 0;
          sin.s <= StartOfFrame;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- start of frame (0xd)
      WHEN StartOfFrame =>
        E_TXD <= x"d";
        E_TX_EN <= '1';

        sin.crc <= x"ffffffff";
        sin.s <= EtherMACDST;

      -- Ethernet DST MAC
      WHEN EtherMACDST =>
        E_TXD <= s.d.dstMAC((s.c * 4 + 3) DOWNTO (s.c * 4));
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(s.d.dstMAC((s.c * 4 + 3) DOWNTO (s.c * 4)), s.crc);
        IF s.c = 11 THEN
          sin.c <= 0;
          sin.s <= EtherMACSRC;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- Ethernet SRC MAC
      WHEN EtherMACSRC =>
        E_TXD <= s.d.srcMAC((s.c * 4 + 3) DOWNTO (s.c * 4));
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(s.d.srcMAC((s.c * 4 + 3) DOWNTO (s.c * 4)), s.crc);
        IF s.c = 11 THEN
          sin.c <= 0;
          sin.s <= EtherType;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- Ethertype 0x0800
      WHEN EtherType =>
        IF s.c = 0 THEN
          E_TXD <= x"8";
          E_TX_EN <= '1';
          sin.crc <= nextCRC32_D4(x"8", s.crc);
          sin.c <= s.c + 1;
        ELSE
          E_TXD <= x"0";
          E_TX_EN <= '1';
          sin.crc <= nextCRC32_D4(x"0", s.crc);
          IF s.c = 3 THEN
            sin.c <= 0;
            sin.s <= IPIHL;
          ELSE
            sin.c <= s.c + 1;
          END IF;
        END IF;

      -- IP IHL 5
      WHEN IPIHL =>
        E_TXD <= x"5";
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(x"5", s.crc);
        sin.c <= 0;
        sin.s <= IPVersion;

      -- IP Version 4
      WHEN IPVersion =>
        E_TXD <= x"4";
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(x"4", s.crc);
        sin.c <= 0;
        sin.s <= IPDSCPECN;

      -- IP DSCP ECN 0x00
      WHEN IPDSCPECN =>
       E_TXD <= x"0";
       E_TX_EN <= '1';
       sin.crc <= nextCRC32_D4(x"0", s.crc);
       IF s.c = 1 THEN
         sin.c <= 0;
         sin.s <= IPLength;
       ELSE
         sin.c <= s.c + 1;
       END IF;

      -- IPLength
      WHEN IPLength =>
        E_TXD <= STD_LOGIC_VECTOR(to_unsigned(s.d.ipLength, E_TXD'length));
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(STD_LOGIC_VECTOR(to_unsigned(s.d.ipLength, E_TXD'length)), s.crc);
        sin.d.ipLength <= s.d.ipLength / 16;
        IF s.c = 3 THEN
          sin.c <= 0;
          sin.s <= IPID;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- IP - ID 0x00
      WHEN IPID =>
        E_TXD <= x"0";
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(x"0", s.crc);
        IF s.c = 3 THEN
          sin.c <= 0;
          sin.s <= IPFlagsFragment;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- IP Flags Fragment Offset 0x00
      WHEN IPFlagsFragment =>
        E_TXD <= x"0";
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(x"0", s.crc);
        IF s.c = 3 THEN
          sin.c <= 0;
          sin.s <= IPTTL;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- IP TTL
      WHEN IPTTL =>
        E_TX_EN <= '1';
        IF s.c = 0 THEN
          E_TXD <= x"0";
          sin.crc <= nextCRC32_D4(x"0", s.crc);
        ELSE
          E_TXD <= x"4";
          sin.crc <= nextCRC32_D4(x"4", s.crc);
        END IF;
        IF s.c = 1 THEN
          sin.c <= 0;
          sin.s <= IPProtocol;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- IP Protocol
      WHEN IPProtocol =>
        E_TXD <= x"1";
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(x"1", s.crc);
        IF s.c = 1 THEN
          sin.c <= 0;
          sin.s <= IPChecksum;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- IPChecksum
      WHEN IPChecksum =>
        E_TXD <= x"0";
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(x"0", s.crc);
        IF s.c = 3 THEN
          sin.c <= 0;
          sin.s <= IPAddrSRC;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- IP Addr SRC
      WHEN IPAddrSRC =>
        E_TXD <= s.d.srcIP((s.c * 4 + 3) DOWNTO (s.c * 4));
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(s.d.srcIP((s.c * 4 + 3) DOWNTO (s.c * 4)), s.crc);
        IF s.c = 7 THEN
          sin.c <= 0;
          sin.s <= IPAddrDST;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- IP Addr DST
      WHEN IPAddrDST =>
        E_TXD <= s.d.dstIP((s.c * 4 + 3) DOWNTO (s.c * 4));
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(s.d.dstIP((s.c * 4 + 3) DOWNTO (s.c * 4)), s.crc);
        IF s.c = 7 THEN
          sin.c <= 0;
          -- Update ME
          sin.s <= DNSMsg;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- UDP Port

      -- DNS Message
      WHEN DNSMsg =>
        E_TXD <= x"C";
        E_TX_EN <= '1';
        sin.crc <= nextCRC32_D4(x"C", s.crc);
        IF s.c = 365 THEN
          sin.c <= 0;
          sin.s <= FrameCheck;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- Ethernet Frame Check Sequence
      WHEN FrameCheck =>
        E_TXD <= NOT s.crc(4 * s.c + 3 DOWNTO 4 * s.c);
        E_TX_EN <= '1';
        IF s.c = 7 THEN
          sin.c <= 0;
          sin.s <= InterframeGap;
        ELSE
          sin.c <= s.c + 1;
        END IF;

      -- Ethernet Interframe Gap
      WHEN InterframeGap =>
        IF s.c = 23 THEN
          sin.c <= 0;
          sin.s <= Idle;
        ELSE
          sin.c <= s.c + 1;
        END IF;
    END CASE;
  END PROCESS;

  snd_reg : PROCESS (E_TX_CLK)
  BEGIN
    IF rising_edge(E_TX_CLK) THEN
      s <= sin;
    END IF;
  END PROCESS;
END rtl;